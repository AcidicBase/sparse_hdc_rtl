// We limit the shift from 1 to 617 (increase later on)
// Note: shift = 0 and shift = HV_DIM are prohibited

// 617 shift values (1 to 617)
parameter integer SHIFTS [0:FEATURE_COUNT-1] = '{247, 51, 125, 429, 478, 113, 299, 545, 283, 100, 453, 446, 4, 112, 407, 
    382, 426, 92, 472, 509, 134, 351, 560, 177, 101, 562, 353, 15, 448, 603, 506, 552, 114, 593, 546, 243, 385, 550, 606, 
    242, 601, 482, 316, 300, 483, 16, 176, 538, 31, 470, 443, 361, 406, 293, 395, 573, 566, 241, 481, 319, 364, 610, 202, 
    592, 62, 43, 1, 501, 223, 273, 37, 126, 12, 305, 473, 78, 72, 47, 567, 508, 544, 17, 88, 217, 197, 240, 33, 454, 557, 
    337, 206, 67, 417, 298, 155, 345, 93, 34, 2, 464, 209, 188, 108, 77, 179, 45, 412, 13, 145, 344, 186, 463, 96, 66, 403, 
    347, 315, 374, 553, 408, 575, 397, 91, 617, 335, 392, 387, 437, 318, 594, 611, 330, 28, 371, 327, 548, 432, 254,198, 
    514, 152, 110, 246, 129, 285, 60, 180, 530, 73, 137, 224, 22, 586, 462, 451, 436, 549, 334, 380, 11, 146, 284, 271,
    466, 457, 280, 411, 372, 389, 433, 516, 439, 350, 504, 409, 477, 87, 38, 118, 488, 50, 230, 294, 303, 500, 604, 35,
    615, 362, 213, 580, 99, 252, 278, 383, 381, 467, 543, 19, 237, 302, 261, 131, 565, 251, 132, 190, 526, 532, 220, 191,
    399, 257, 450, 68, 613, 75, 235, 227, 222, 554, 355, 154, 57, 279, 400, 542, 484, 103, 491, 311, 116, 533, 249, 605, 
    324, 297, 104, 30, 596, 123, 569, 168, 313, 162, 499, 258, 83, 74, 182, 140, 614, 270, 321, 158, 591, 189, 358, 430, 
    183, 486, 82, 42, 232, 348, 394, 26, 54, 578, 519, 539, 151, 495, 398, 195, 63, 431, 317, 413, 304, 590, 205, 124, 521, 
    352, 218, 55, 141, 120, 338, 584, 178, 208, 262, 375, 153, 474, 328, 27, 89, 365, 6, 65, 607, 452, 185, 58, 515, 139, 
    250, 225, 21, 292, 609, 76, 354, 289, 90, 111, 494, 568, 107, 363, 574, 422, 511, 143, 40, 119, 558, 290, 256, 69, 551, 
    570, 536, 600, 253, 410, 277, 268, 428, 48, 18, 266, 64, 25, 359, 518, 421, 142, 39, 336, 148, 231, 534, 458, 420, 115, 
    7, 296, 340, 32, 117, 333, 135, 404, 331, 10, 465, 479, 163, 309, 80, 204, 447, 563, 173, 286, 147, 555, 487, 571, 438, 
    171, 349, 440, 71, 390, 459, 480, 402, 391, 329, 384, 377, 595, 200, 194, 524, 128, 424, 489, 275, 23, 416, 492, 36, 556, 
    84, 517, 3, 184, 370, 540, 207, 150, 496, 144, 79, 109, 577, 199, 105, 248, 396, 267, 165, 5, 427, 561, 226, 461, 388, 
    234, 136, 612, 341, 493, 378, 513, 525, 583, 582, 520, 215, 547, 122, 343, 598, 260, 523, 528, 174, 212, 169, 423, 167, 
    20, 216, 201, 356, 81, 323, 44, 367, 531, 444, 228, 9, 265, 326, 8, 86, 70, 166, 342, 170, 274, 322, 59, 449, 203, 157, 
    181, 376, 221, 469, 527, 587, 339, 597, 192, 127, 535, 29, 98, 160, 386, 507, 456, 346, 53, 541, 608, 485, 442, 441, 244, 
    529, 476, 133, 585, 366, 360, 581, 56, 589, 196, 161, 85, 471, 156, 502, 616, 95, 172, 295, 263, 312, 320, 576, 435, 405, 
    497, 559, 210, 425, 368, 106, 434, 579, 264, 415, 159, 238, 236, 588, 149, 269, 307, 61, 130, 325, 164, 288, 41, 193, 233, 
    418, 245, 455, 393, 314, 282, 49, 97, 276, 46, 503, 102, 175, 572, 94, 229, 602, 219, 445, 310, 369, 505, 510, 522, 498, 
    490, 537, 255, 460, 52, 272, 239, 259, 373, 287, 281, 308, 211, 187, 332, 301, 121, 24, 512, 401, 291, 357, 475, 419, 14, 
    468, 564, 414, 379, 599, 214, 138, 306}; 
