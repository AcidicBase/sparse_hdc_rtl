module IM_Output_Switch(output_id, level_hv, input_hv);
  input [3:0] output_id;
  input [9:0] output_hv;
  output reg [616:0][9:0] level_hv;

  always@(*) begin
    case(output_id)
      0 : level_hv[0][9:0] = output_hv;
      1 : level_hv[1][9:0] = output_hv;
      2 : level_hv[2][9:0] = output_hv;
      3 : level_hv[3][9:0] = output_hv;
      4 : level_hv[4][9:0] = output_hv;
      5 : level_hv[5][9:0] = output_hv;
      6 : level_hv[6][9:0] = output_hv;
      7 : level_hv[7][9:0] = output_hv;
      8 : level_hv[8][9:0] = output_hv;
      9 : level_hv[9][9:0] = output_hv;
      10 : level_hv[10][9:0] = output_hv;
      11 : level_hv[11][9:0] = output_hv;
      12 : level_hv[12][9:0] = output_hv;
      13 : level_hv[13][9:0] = output_hv;
      14 : level_hv[14][9:0] = output_hv;
      15 : level_hv[15][9:0] = output_hv;
      16 : level_hv[16][9:0] = output_hv;
      17 : level_hv[17][9:0] = output_hv;
      18 : level_hv[18][9:0] = output_hv;
      19 : level_hv[19][9:0] = output_hv;
      20 : level_hv[20][9:0] = output_hv;
      21 : level_hv[21][9:0] = output_hv;
      22 : level_hv[22][9:0] = output_hv;
      23 : level_hv[23][9:0] = output_hv;
      24 : level_hv[24][9:0] = output_hv;
      25 : level_hv[25][9:0] = output_hv;
      26 : level_hv[26][9:0] = output_hv;
      27 : level_hv[27][9:0] = output_hv;
      28 : level_hv[28][9:0] = output_hv;
      29 : level_hv[29][9:0] = output_hv;
      30 : level_hv[30][9:0] = output_hv;
      31 : level_hv[31][9:0] = output_hv;
      32 : level_hv[32][9:0] = output_hv;
      33 : level_hv[33][9:0] = output_hv;
      34 : level_hv[34][9:0] = output_hv;
      35 : level_hv[35][9:0] = output_hv;
      36 : level_hv[36][9:0] = output_hv;
      37 : level_hv[37][9:0] = output_hv;
      38 : level_hv[38][9:0] = output_hv;
      39 : level_hv[39][9:0] = output_hv;
      40 : level_hv[40][9:0] = output_hv;
      41 : level_hv[41][9:0] = output_hv;
      42 : level_hv[42][9:0] = output_hv;
      43 : level_hv[43][9:0] = output_hv;
      44 : level_hv[44][9:0] = output_hv;
      45 : level_hv[45][9:0] = output_hv;
      46 : level_hv[46][9:0] = output_hv;
      47 : level_hv[47][9:0] = output_hv;
      48 : level_hv[48][9:0] = output_hv;
      49 : level_hv[49][9:0] = output_hv;
      50 : level_hv[50][9:0] = output_hv;
      51 : level_hv[51][9:0] = output_hv;
      52 : level_hv[52][9:0] = output_hv;
      53 : level_hv[53][9:0] = output_hv;
      54 : level_hv[54][9:0] = output_hv;
      55 : level_hv[55][9:0] = output_hv;
      56 : level_hv[56][9:0] = output_hv;
      57 : level_hv[57][9:0] = output_hv;
      58 : level_hv[58][9:0] = output_hv;
      59 : level_hv[59][9:0] = output_hv;
      60 : level_hv[60][9:0] = output_hv;
      61 : level_hv[61][9:0] = output_hv;
      62 : level_hv[62][9:0] = output_hv;
      63 : level_hv[63][9:0] = output_hv;
      64 : level_hv[64][9:0] = output_hv;
      65 : level_hv[65][9:0] = output_hv;
      66 : level_hv[66][9:0] = output_hv;
      67 : level_hv[67][9:0] = output_hv;
      68 : level_hv[68][9:0] = output_hv;
      69 : level_hv[69][9:0] = output_hv;
      70 : level_hv[70][9:0] = output_hv;
      71 : level_hv[71][9:0] = output_hv;
      72 : level_hv[72][9:0] = output_hv;
      73 : level_hv[73][9:0] = output_hv;
      74 : level_hv[74][9:0] = output_hv;
      75 : level_hv[75][9:0] = output_hv;
      76 : level_hv[76][9:0] = output_hv;
      77 : level_hv[77][9:0] = output_hv;
      78 : level_hv[78][9:0] = output_hv;
      79 : level_hv[79][9:0] = output_hv;
      80 : level_hv[80][9:0] = output_hv;
      81 : level_hv[81][9:0] = output_hv;
      82 : level_hv[82][9:0] = output_hv;
      83 : level_hv[83][9:0] = output_hv;
      84 : level_hv[84][9:0] = output_hv;
      85 : level_hv[85][9:0] = output_hv;
      86 : level_hv[86][9:0] = output_hv;
      87 : level_hv[87][9:0] = output_hv;
      88 : level_hv[88][9:0] = output_hv;
      89 : level_hv[89][9:0] = output_hv;
      90 : level_hv[90][9:0] = output_hv;
      91 : level_hv[91][9:0] = output_hv;
      92 : level_hv[92][9:0] = output_hv;
      93 : level_hv[93][9:0] = output_hv;
      94 : level_hv[94][9:0] = output_hv;
      95 : level_hv[95][9:0] = output_hv;
      96 : level_hv[96][9:0] = output_hv;
      97 : level_hv[97][9:0] = output_hv;
      98 : level_hv[98][9:0] = output_hv;
      99 : level_hv[99][9:0] = output_hv;
      100 : level_hv[100][9:0] = output_hv;
      101 : level_hv[101][9:0] = output_hv;
      102 : level_hv[102][9:0] = output_hv;
      103 : level_hv[103][9:0] = output_hv;
      104 : level_hv[104][9:0] = output_hv;
      105 : level_hv[105][9:0] = output_hv;
      106 : level_hv[106][9:0] = output_hv;
      107 : level_hv[107][9:0] = output_hv;
      108 : level_hv[108][9:0] = output_hv;
      109 : level_hv[109][9:0] = output_hv;
      110 : level_hv[110][9:0] = output_hv;
      111 : level_hv[111][9:0] = output_hv;
      112 : level_hv[112][9:0] = output_hv;
      113 : level_hv[113][9:0] = output_hv;
      114 : level_hv[114][9:0] = output_hv;
      115 : level_hv[115][9:0] = output_hv;
      116 : level_hv[116][9:0] = output_hv;
      117 : level_hv[117][9:0] = output_hv;
      118 : level_hv[118][9:0] = output_hv;
      119 : level_hv[119][9:0] = output_hv;
      120 : level_hv[120][9:0] = output_hv;
      121 : level_hv[121][9:0] = output_hv;
      122 : level_hv[122][9:0] = output_hv;
      123 : level_hv[123][9:0] = output_hv;
      124 : level_hv[124][9:0] = output_hv;
      125 : level_hv[125][9:0] = output_hv;
      126 : level_hv[126][9:0] = output_hv;
      127 : level_hv[127][9:0] = output_hv;
      128 : level_hv[128][9:0] = output_hv;
      129 : level_hv[129][9:0] = output_hv;
      130 : level_hv[130][9:0] = output_hv;
      131 : level_hv[131][9:0] = output_hv;
      132 : level_hv[132][9:0] = output_hv;
      133 : level_hv[133][9:0] = output_hv;
      134 : level_hv[134][9:0] = output_hv;
      135 : level_hv[135][9:0] = output_hv;
      136 : level_hv[136][9:0] = output_hv;
      137 : level_hv[137][9:0] = output_hv;
      138 : level_hv[138][9:0] = output_hv;
      139 : level_hv[139][9:0] = output_hv;
      140 : level_hv[140][9:0] = output_hv;
      141 : level_hv[141][9:0] = output_hv;
      142 : level_hv[142][9:0] = output_hv;
      143 : level_hv[143][9:0] = output_hv;
      144 : level_hv[144][9:0] = output_hv;
      145 : level_hv[145][9:0] = output_hv;
      146 : level_hv[146][9:0] = output_hv;
      147 : level_hv[147][9:0] = output_hv;
      148 : level_hv[148][9:0] = output_hv;
      149 : level_hv[149][9:0] = output_hv;
      150 : level_hv[150][9:0] = output_hv;
      151 : level_hv[151][9:0] = output_hv;
      152 : level_hv[152][9:0] = output_hv;
      153 : level_hv[153][9:0] = output_hv;
      154 : level_hv[154][9:0] = output_hv;
      155 : level_hv[155][9:0] = output_hv;
      156 : level_hv[156][9:0] = output_hv;
      157 : level_hv[157][9:0] = output_hv;
      158 : level_hv[158][9:0] = output_hv;
      159 : level_hv[159][9:0] = output_hv;
      160 : level_hv[160][9:0] = output_hv;
      161 : level_hv[161][9:0] = output_hv;
      162 : level_hv[162][9:0] = output_hv;
      163 : level_hv[163][9:0] = output_hv;
      164 : level_hv[164][9:0] = output_hv;
      165 : level_hv[165][9:0] = output_hv;
      166 : level_hv[166][9:0] = output_hv;
      167 : level_hv[167][9:0] = output_hv;
      168 : level_hv[168][9:0] = output_hv;
      169 : level_hv[169][9:0] = output_hv;
      170 : level_hv[170][9:0] = output_hv;
      171 : level_hv[171][9:0] = output_hv;
      172 : level_hv[172][9:0] = output_hv;
      173 : level_hv[173][9:0] = output_hv;
      174 : level_hv[174][9:0] = output_hv;
      175 : level_hv[175][9:0] = output_hv;
      176 : level_hv[176][9:0] = output_hv;
      177 : level_hv[177][9:0] = output_hv;
      178 : level_hv[178][9:0] = output_hv;
      179 : level_hv[179][9:0] = output_hv;
      180 : level_hv[180][9:0] = output_hv;
      181 : level_hv[181][9:0] = output_hv;
      182 : level_hv[182][9:0] = output_hv;
      183 : level_hv[183][9:0] = output_hv;
      184 : level_hv[184][9:0] = output_hv;
      185 : level_hv[185][9:0] = output_hv;
      186 : level_hv[186][9:0] = output_hv;
      187 : level_hv[187][9:0] = output_hv;
      188 : level_hv[188][9:0] = output_hv;
      189 : level_hv[189][9:0] = output_hv;
      190 : level_hv[190][9:0] = output_hv;
      191 : level_hv[191][9:0] = output_hv;
      192 : level_hv[192][9:0] = output_hv;
      193 : level_hv[193][9:0] = output_hv;
      194 : level_hv[194][9:0] = output_hv;
      195 : level_hv[195][9:0] = output_hv;
      196 : level_hv[196][9:0] = output_hv;
      197 : level_hv[197][9:0] = output_hv;
      198 : level_hv[198][9:0] = output_hv;
      199 : level_hv[199][9:0] = output_hv;
      200 : level_hv[200][9:0] = output_hv;
      201 : level_hv[201][9:0] = output_hv;
      202 : level_hv[202][9:0] = output_hv;
      203 : level_hv[203][9:0] = output_hv;
      204 : level_hv[204][9:0] = output_hv;
      205 : level_hv[205][9:0] = output_hv;
      206 : level_hv[206][9:0] = output_hv;
      207 : level_hv[207][9:0] = output_hv;
      208 : level_hv[208][9:0] = output_hv;
      209 : level_hv[209][9:0] = output_hv;
      210 : level_hv[210][9:0] = output_hv;
      211 : level_hv[211][9:0] = output_hv;
      212 : level_hv[212][9:0] = output_hv;
      213 : level_hv[213][9:0] = output_hv;
      214 : level_hv[214][9:0] = output_hv;
      215 : level_hv[215][9:0] = output_hv;
      216 : level_hv[216][9:0] = output_hv;
      217 : level_hv[217][9:0] = output_hv;
      218 : level_hv[218][9:0] = output_hv;
      219 : level_hv[219][9:0] = output_hv;
      220 : level_hv[220][9:0] = output_hv;
      221 : level_hv[221][9:0] = output_hv;
      222 : level_hv[222][9:0] = output_hv;
      223 : level_hv[223][9:0] = output_hv;
      224 : level_hv[224][9:0] = output_hv;
      225 : level_hv[225][9:0] = output_hv;
      226 : level_hv[226][9:0] = output_hv;
      227 : level_hv[227][9:0] = output_hv;
      228 : level_hv[228][9:0] = output_hv;
      229 : level_hv[229][9:0] = output_hv;
      230 : level_hv[230][9:0] = output_hv;
      231 : level_hv[231][9:0] = output_hv;
      232 : level_hv[232][9:0] = output_hv;
      233 : level_hv[233][9:0] = output_hv;
      234 : level_hv[234][9:0] = output_hv;
      235 : level_hv[235][9:0] = output_hv;
      236 : level_hv[236][9:0] = output_hv;
      237 : level_hv[237][9:0] = output_hv;
      238 : level_hv[238][9:0] = output_hv;
      239 : level_hv[239][9:0] = output_hv;
      240 : level_hv[240][9:0] = output_hv;
      241 : level_hv[241][9:0] = output_hv;
      242 : level_hv[242][9:0] = output_hv;
      243 : level_hv[243][9:0] = output_hv;
      244 : level_hv[244][9:0] = output_hv;
      245 : level_hv[245][9:0] = output_hv;
      246 : level_hv[246][9:0] = output_hv;
      247 : level_hv[247][9:0] = output_hv;
      248 : level_hv[248][9:0] = output_hv;
      249 : level_hv[249][9:0] = output_hv;
      250 : level_hv[250][9:0] = output_hv;
      251 : level_hv[251][9:0] = output_hv;
      252 : level_hv[252][9:0] = output_hv;
      253 : level_hv[253][9:0] = output_hv;
      254 : level_hv[254][9:0] = output_hv;
      255 : level_hv[255][9:0] = output_hv;
      256 : level_hv[256][9:0] = output_hv;
      257 : level_hv[257][9:0] = output_hv;
      258 : level_hv[258][9:0] = output_hv;
      259 : level_hv[259][9:0] = output_hv;
      260 : level_hv[260][9:0] = output_hv;
      261 : level_hv[261][9:0] = output_hv;
      262 : level_hv[262][9:0] = output_hv;
      263 : level_hv[263][9:0] = output_hv;
      264 : level_hv[264][9:0] = output_hv;
      265 : level_hv[265][9:0] = output_hv;
      266 : level_hv[266][9:0] = output_hv;
      267 : level_hv[267][9:0] = output_hv;
      268 : level_hv[268][9:0] = output_hv;
      269 : level_hv[269][9:0] = output_hv;
      270 : level_hv[270][9:0] = output_hv;
      271 : level_hv[271][9:0] = output_hv;
      272 : level_hv[272][9:0] = output_hv;
      273 : level_hv[273][9:0] = output_hv;
      274 : level_hv[274][9:0] = output_hv;
      275 : level_hv[275][9:0] = output_hv;
      276 : level_hv[276][9:0] = output_hv;
      277 : level_hv[277][9:0] = output_hv;
      278 : level_hv[278][9:0] = output_hv;
      279 : level_hv[279][9:0] = output_hv;
      280 : level_hv[280][9:0] = output_hv;
      281 : level_hv[281][9:0] = output_hv;
      282 : level_hv[282][9:0] = output_hv;
      283 : level_hv[283][9:0] = output_hv;
      284 : level_hv[284][9:0] = output_hv;
      285 : level_hv[285][9:0] = output_hv;
      286 : level_hv[286][9:0] = output_hv;
      287 : level_hv[287][9:0] = output_hv;
      288 : level_hv[288][9:0] = output_hv;
      289 : level_hv[289][9:0] = output_hv;
      290 : level_hv[290][9:0] = output_hv;
      291 : level_hv[291][9:0] = output_hv;
      292 : level_hv[292][9:0] = output_hv;
      293 : level_hv[293][9:0] = output_hv;
      294 : level_hv[294][9:0] = output_hv;
      295 : level_hv[295][9:0] = output_hv;
      296 : level_hv[296][9:0] = output_hv;
      297 : level_hv[297][9:0] = output_hv;
      298 : level_hv[298][9:0] = output_hv;
      299 : level_hv[299][9:0] = output_hv;
      300 : level_hv[300][9:0] = output_hv;
      301 : level_hv[301][9:0] = output_hv;
      302 : level_hv[302][9:0] = output_hv;
      303 : level_hv[303][9:0] = output_hv;
      304 : level_hv[304][9:0] = output_hv;
      305 : level_hv[305][9:0] = output_hv;
      306 : level_hv[306][9:0] = output_hv;
      307 : level_hv[307][9:0] = output_hv;
      308 : level_hv[308][9:0] = output_hv;
      309 : level_hv[309][9:0] = output_hv;
      310 : level_hv[310][9:0] = output_hv;
      311 : level_hv[311][9:0] = output_hv;
      312 : level_hv[312][9:0] = output_hv;
      313 : level_hv[313][9:0] = output_hv;
      314 : level_hv[314][9:0] = output_hv;
      315 : level_hv[315][9:0] = output_hv;
      316 : level_hv[316][9:0] = output_hv;
      317 : level_hv[317][9:0] = output_hv;
      318 : level_hv[318][9:0] = output_hv;
      319 : level_hv[319][9:0] = output_hv;
      320 : level_hv[320][9:0] = output_hv;
      321 : level_hv[321][9:0] = output_hv;
      322 : level_hv[322][9:0] = output_hv;
      323 : level_hv[323][9:0] = output_hv;
      324 : level_hv[324][9:0] = output_hv;
      325 : level_hv[325][9:0] = output_hv;
      326 : level_hv[326][9:0] = output_hv;
      327 : level_hv[327][9:0] = output_hv;
      328 : level_hv[328][9:0] = output_hv;
      329 : level_hv[329][9:0] = output_hv;
      330 : level_hv[330][9:0] = output_hv;
      331 : level_hv[331][9:0] = output_hv;
      332 : level_hv[332][9:0] = output_hv;
      333 : level_hv[333][9:0] = output_hv;
      334 : level_hv[334][9:0] = output_hv;
      335 : level_hv[335][9:0] = output_hv;
      336 : level_hv[336][9:0] = output_hv;
      337 : level_hv[337][9:0] = output_hv;
      338 : level_hv[338][9:0] = output_hv;
      339 : level_hv[339][9:0] = output_hv;
      340 : level_hv[340][9:0] = output_hv;
      341 : level_hv[341][9:0] = output_hv;
      342 : level_hv[342][9:0] = output_hv;
      343 : level_hv[343][9:0] = output_hv;
      344 : level_hv[344][9:0] = output_hv;
      345 : level_hv[345][9:0] = output_hv;
      346 : level_hv[346][9:0] = output_hv;
      347 : level_hv[347][9:0] = output_hv;
      348 : level_hv[348][9:0] = output_hv;
      349 : level_hv[349][9:0] = output_hv;
      350 : level_hv[350][9:0] = output_hv;
      351 : level_hv[351][9:0] = output_hv;
      352 : level_hv[352][9:0] = output_hv;
      353 : level_hv[353][9:0] = output_hv;
      354 : level_hv[354][9:0] = output_hv;
      355 : level_hv[355][9:0] = output_hv;
      356 : level_hv[356][9:0] = output_hv;
      357 : level_hv[357][9:0] = output_hv;
      358 : level_hv[358][9:0] = output_hv;
      359 : level_hv[359][9:0] = output_hv;
      360 : level_hv[360][9:0] = output_hv;
      361 : level_hv[361][9:0] = output_hv;
      362 : level_hv[362][9:0] = output_hv;
      363 : level_hv[363][9:0] = output_hv;
      364 : level_hv[364][9:0] = output_hv;
      365 : level_hv[365][9:0] = output_hv;
      366 : level_hv[366][9:0] = output_hv;
      367 : level_hv[367][9:0] = output_hv;
      368 : level_hv[368][9:0] = output_hv;
      369 : level_hv[369][9:0] = output_hv;
      370 : level_hv[370][9:0] = output_hv;
      371 : level_hv[371][9:0] = output_hv;
      372 : level_hv[372][9:0] = output_hv;
      373 : level_hv[373][9:0] = output_hv;
      374 : level_hv[374][9:0] = output_hv;
      375 : level_hv[375][9:0] = output_hv;
      376 : level_hv[376][9:0] = output_hv;
      377 : level_hv[377][9:0] = output_hv;
      378 : level_hv[378][9:0] = output_hv;
      379 : level_hv[379][9:0] = output_hv;
      380 : level_hv[380][9:0] = output_hv;
      381 : level_hv[381][9:0] = output_hv;
      382 : level_hv[382][9:0] = output_hv;
      383 : level_hv[383][9:0] = output_hv;
      384 : level_hv[384][9:0] = output_hv;
      385 : level_hv[385][9:0] = output_hv;
      386 : level_hv[386][9:0] = output_hv;
      387 : level_hv[387][9:0] = output_hv;
      388 : level_hv[388][9:0] = output_hv;
      389 : level_hv[389][9:0] = output_hv;
      390 : level_hv[390][9:0] = output_hv;
      391 : level_hv[391][9:0] = output_hv;
      392 : level_hv[392][9:0] = output_hv;
      393 : level_hv[393][9:0] = output_hv;
      394 : level_hv[394][9:0] = output_hv;
      395 : level_hv[395][9:0] = output_hv;
      396 : level_hv[396][9:0] = output_hv;
      397 : level_hv[397][9:0] = output_hv;
      398 : level_hv[398][9:0] = output_hv;
      399 : level_hv[399][9:0] = output_hv;
      400 : level_hv[400][9:0] = output_hv;
      401 : level_hv[401][9:0] = output_hv;
      402 : level_hv[402][9:0] = output_hv;
      403 : level_hv[403][9:0] = output_hv;
      404 : level_hv[404][9:0] = output_hv;
      405 : level_hv[405][9:0] = output_hv;
      406 : level_hv[406][9:0] = output_hv;
      407 : level_hv[407][9:0] = output_hv;
      408 : level_hv[408][9:0] = output_hv;
      409 : level_hv[409][9:0] = output_hv;
      410 : level_hv[410][9:0] = output_hv;
      411 : level_hv[411][9:0] = output_hv;
      412 : level_hv[412][9:0] = output_hv;
      413 : level_hv[413][9:0] = output_hv;
      414 : level_hv[414][9:0] = output_hv;
      415 : level_hv[415][9:0] = output_hv;
      416 : level_hv[416][9:0] = output_hv;
      417 : level_hv[417][9:0] = output_hv;
      418 : level_hv[418][9:0] = output_hv;
      419 : level_hv[419][9:0] = output_hv;
      420 : level_hv[420][9:0] = output_hv;
      421 : level_hv[421][9:0] = output_hv;
      422 : level_hv[422][9:0] = output_hv;
      423 : level_hv[423][9:0] = output_hv;
      424 : level_hv[424][9:0] = output_hv;
      425 : level_hv[425][9:0] = output_hv;
      426 : level_hv[426][9:0] = output_hv;
      427 : level_hv[427][9:0] = output_hv;
      428 : level_hv[428][9:0] = output_hv;
      429 : level_hv[429][9:0] = output_hv;
      430 : level_hv[430][9:0] = output_hv;
      431 : level_hv[431][9:0] = output_hv;
      432 : level_hv[432][9:0] = output_hv;
      433 : level_hv[433][9:0] = output_hv;
      434 : level_hv[434][9:0] = output_hv;
      435 : level_hv[435][9:0] = output_hv;
      436 : level_hv[436][9:0] = output_hv;
      437 : level_hv[437][9:0] = output_hv;
      438 : level_hv[438][9:0] = output_hv;
      439 : level_hv[439][9:0] = output_hv;
      440 : level_hv[440][9:0] = output_hv;
      441 : level_hv[441][9:0] = output_hv;
      442 : level_hv[442][9:0] = output_hv;
      443 : level_hv[443][9:0] = output_hv;
      444 : level_hv[444][9:0] = output_hv;
      445 : level_hv[445][9:0] = output_hv;
      446 : level_hv[446][9:0] = output_hv;
      447 : level_hv[447][9:0] = output_hv;
      448 : level_hv[448][9:0] = output_hv;
      449 : level_hv[449][9:0] = output_hv;
      450 : level_hv[450][9:0] = output_hv;
      451 : level_hv[451][9:0] = output_hv;
      452 : level_hv[452][9:0] = output_hv;
      453 : level_hv[453][9:0] = output_hv;
      454 : level_hv[454][9:0] = output_hv;
      455 : level_hv[455][9:0] = output_hv;
      456 : level_hv[456][9:0] = output_hv;
      457 : level_hv[457][9:0] = output_hv;
      458 : level_hv[458][9:0] = output_hv;
      459 : level_hv[459][9:0] = output_hv;
      460 : level_hv[460][9:0] = output_hv;
      461 : level_hv[461][9:0] = output_hv;
      462 : level_hv[462][9:0] = output_hv;
      463 : level_hv[463][9:0] = output_hv;
      464 : level_hv[464][9:0] = output_hv;
      465 : level_hv[465][9:0] = output_hv;
      466 : level_hv[466][9:0] = output_hv;
      467 : level_hv[467][9:0] = output_hv;
      468 : level_hv[468][9:0] = output_hv;
      469 : level_hv[469][9:0] = output_hv;
      470 : level_hv[470][9:0] = output_hv;
      471 : level_hv[471][9:0] = output_hv;
      472 : level_hv[472][9:0] = output_hv;
      473 : level_hv[473][9:0] = output_hv;
      474 : level_hv[474][9:0] = output_hv;
      475 : level_hv[475][9:0] = output_hv;
      476 : level_hv[476][9:0] = output_hv;
      477 : level_hv[477][9:0] = output_hv;
      478 : level_hv[478][9:0] = output_hv;
      479 : level_hv[479][9:0] = output_hv;
      480 : level_hv[480][9:0] = output_hv;
      481 : level_hv[481][9:0] = output_hv;
      482 : level_hv[482][9:0] = output_hv;
      483 : level_hv[483][9:0] = output_hv;
      484 : level_hv[484][9:0] = output_hv;
      485 : level_hv[485][9:0] = output_hv;
      486 : level_hv[486][9:0] = output_hv;
      487 : level_hv[487][9:0] = output_hv;
      488 : level_hv[488][9:0] = output_hv;
      489 : level_hv[489][9:0] = output_hv;
      490 : level_hv[490][9:0] = output_hv;
      491 : level_hv[491][9:0] = output_hv;
      492 : level_hv[492][9:0] = output_hv;
      493 : level_hv[493][9:0] = output_hv;
      494 : level_hv[494][9:0] = output_hv;
      495 : level_hv[495][9:0] = output_hv;
      496 : level_hv[496][9:0] = output_hv;
      497 : level_hv[497][9:0] = output_hv;
      498 : level_hv[498][9:0] = output_hv;
      499 : level_hv[499][9:0] = output_hv;
      500 : level_hv[500][9:0] = output_hv;
      501 : level_hv[501][9:0] = output_hv;
      502 : level_hv[502][9:0] = output_hv;
      503 : level_hv[503][9:0] = output_hv;
      504 : level_hv[504][9:0] = output_hv;
      505 : level_hv[505][9:0] = output_hv;
      506 : level_hv[506][9:0] = output_hv;
      507 : level_hv[507][9:0] = output_hv;
      508 : level_hv[508][9:0] = output_hv;
      509 : level_hv[509][9:0] = output_hv;
      510 : level_hv[510][9:0] = output_hv;
      511 : level_hv[511][9:0] = output_hv;
      512 : level_hv[512][9:0] = output_hv;
      513 : level_hv[513][9:0] = output_hv;
      514 : level_hv[514][9:0] = output_hv;
      515 : level_hv[515][9:0] = output_hv;
      516 : level_hv[516][9:0] = output_hv;
      517 : level_hv[517][9:0] = output_hv;
      518 : level_hv[518][9:0] = output_hv;
      519 : level_hv[519][9:0] = output_hv;
      520 : level_hv[520][9:0] = output_hv;
      521 : level_hv[521][9:0] = output_hv;
      522 : level_hv[522][9:0] = output_hv;
      523 : level_hv[523][9:0] = output_hv;
      524 : level_hv[524][9:0] = output_hv;
      525 : level_hv[525][9:0] = output_hv;
      526 : level_hv[526][9:0] = output_hv;
      527 : level_hv[527][9:0] = output_hv;
      528 : level_hv[528][9:0] = output_hv;
      529 : level_hv[529][9:0] = output_hv;
      530 : level_hv[530][9:0] = output_hv;
      531 : level_hv[531][9:0] = output_hv;
      532 : level_hv[532][9:0] = output_hv;
      533 : level_hv[533][9:0] = output_hv;
      534 : level_hv[534][9:0] = output_hv;
      535 : level_hv[535][9:0] = output_hv;
      536 : level_hv[536][9:0] = output_hv;
      537 : level_hv[537][9:0] = output_hv;
      538 : level_hv[538][9:0] = output_hv;
      539 : level_hv[539][9:0] = output_hv;
      540 : level_hv[540][9:0] = output_hv;
      541 : level_hv[541][9:0] = output_hv;
      542 : level_hv[542][9:0] = output_hv;
      543 : level_hv[543][9:0] = output_hv;
      544 : level_hv[544][9:0] = output_hv;
      545 : level_hv[545][9:0] = output_hv;
      546 : level_hv[546][9:0] = output_hv;
      547 : level_hv[547][9:0] = output_hv;
      548 : level_hv[548][9:0] = output_hv;
      549 : level_hv[549][9:0] = output_hv;
      550 : level_hv[550][9:0] = output_hv;
      551 : level_hv[551][9:0] = output_hv;
      552 : level_hv[552][9:0] = output_hv;
      553 : level_hv[553][9:0] = output_hv;
      554 : level_hv[554][9:0] = output_hv;
      555 : level_hv[555][9:0] = output_hv;
      556 : level_hv[556][9:0] = output_hv;
      557 : level_hv[557][9:0] = output_hv;
      558 : level_hv[558][9:0] = output_hv;
      559 : level_hv[559][9:0] = output_hv;
      560 : level_hv[560][9:0] = output_hv;
      561 : level_hv[561][9:0] = output_hv;
      562 : level_hv[562][9:0] = output_hv;
      563 : level_hv[563][9:0] = output_hv;
      564 : level_hv[564][9:0] = output_hv;
      565 : level_hv[565][9:0] = output_hv;
      566 : level_hv[566][9:0] = output_hv;
      567 : level_hv[567][9:0] = output_hv;
      568 : level_hv[568][9:0] = output_hv;
      569 : level_hv[569][9:0] = output_hv;
      570 : level_hv[570][9:0] = output_hv;
      571 : level_hv[571][9:0] = output_hv;
      572 : level_hv[572][9:0] = output_hv;
      573 : level_hv[573][9:0] = output_hv;
      574 : level_hv[574][9:0] = output_hv;
      575 : level_hv[575][9:0] = output_hv;
      576 : level_hv[576][9:0] = output_hv;
      577 : level_hv[577][9:0] = output_hv;
      578 : level_hv[578][9:0] = output_hv;
      579 : level_hv[579][9:0] = output_hv;
      580 : level_hv[580][9:0] = output_hv;
      581 : level_hv[581][9:0] = output_hv;
      582 : level_hv[582][9:0] = output_hv;
      583 : level_hv[583][9:0] = output_hv;
      584 : level_hv[584][9:0] = output_hv;
      585 : level_hv[585][9:0] = output_hv;
      586 : level_hv[586][9:0] = output_hv;
      587 : level_hv[587][9:0] = output_hv;
      588 : level_hv[588][9:0] = output_hv;
      589 : level_hv[589][9:0] = output_hv;
      590 : level_hv[590][9:0] = output_hv;
      591 : level_hv[591][9:0] = output_hv;
      592 : level_hv[592][9:0] = output_hv;
      593 : level_hv[593][9:0] = output_hv;
      594 : level_hv[594][9:0] = output_hv;
      595 : level_hv[595][9:0] = output_hv;
      596 : level_hv[596][9:0] = output_hv;
      597 : level_hv[597][9:0] = output_hv;
      598 : level_hv[598][9:0] = output_hv;
      599 : level_hv[599][9:0] = output_hv;
      600 : level_hv[600][9:0] = output_hv;
      601 : level_hv[601][9:0] = output_hv;
      602 : level_hv[602][9:0] = output_hv;
      603 : level_hv[603][9:0] = output_hv;
      604 : level_hv[604][9:0] = output_hv;
      605 : level_hv[605][9:0] = output_hv;
      606 : level_hv[606][9:0] = output_hv;
      607 : level_hv[607][9:0] = output_hv;
      608 : level_hv[608][9:0] = output_hv;
      609 : level_hv[609][9:0] = output_hv;
      610 : level_hv[610][9:0] = output_hv;
      611 : level_hv[611][9:0] = output_hv;
      612 : level_hv[612][9:0] = output_hv;
      613 : level_hv[613][9:0] = output_hv;
      614 : level_hv[614][9:0] = output_hv;
      615 : level_hv[615][9:0] = output_hv;
      616 : level_hv[616][9:0] = output_hv;
    endcase
  end
endmodule

