// `include "TB_Quantizer.sv"
// `include "TB_FLOAT32_Comparator.sv"
// `include "TB_IM_Fetch.sv"
`include "TB_Encoder.sv"