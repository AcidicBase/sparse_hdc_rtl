`timescale 1ns / 1ps

module assoc_tree_adder(

    );
endmodule
